// Contains the immediate parameters for the immediate generation unit of RISC-V RS32IM

`ifndef IMMPARAMETERS_VH
`define IMMPARAMETERS_VH

// Immediate parameters
`define ITypeImm 2'b00
`define STypeImm 2'b01
`define UTypeImm 2'b10

`endif